// And Gate
module and_gate(
	input wire a, b,
	output wire c
	);
	assign c = a & b;
endmodule
